----------------------------------------------------------------------------------
-- Engineer: Mike Field <hamster@snap.net.nz>
-- 
-- Description: Generate analog 800x600 VGA, double-doublescanned from 19200 bytes of RAM
--
-- see http://hamsterworks.co.nz/mediawiki/index.php/OV7670_camera for more information
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity vga_disp is
    Port ( 
      clk50       : in  STD_LOGIC;
	  vga_state	  : in  STD_LOGIC;
	  vga_shift	  : in  STD_LOGIC;
      vga_red     : out STD_LOGIC;
      vga_green   : out STD_LOGIC;
      vga_blue    : out STD_LOGIC;
      vga_hsync   : out STD_LOGIC;
      vga_vsync   : out STD_LOGIC
    );
end vga_disp;

architecture Behavioral of vga_disp is
   -- Timing constants
   constant hRez       : natural := 800;
   constant vRez       : natural := 600;

   constant hMaxCount  : natural := 1056;
   constant hStartSync : natural := 928;
   constant hEndSync   : natural := 1056;
   constant vMaxCount  : natural := 628;
   constant vStartSync : natural := 624;
   constant vEndSync   : natural := 628;
   constant hsync_active : std_logic := '0';
   constant vsync_active : std_logic := '0';

   signal hCounter : unsigned(10 downto 0) := (others => '0');
   signal vCounter : unsigned(9 downto 0) := (others => '0');
   signal hdispCounter : unsigned(2 downto 0) := (others => '0');
   signal vdispCounter : unsigned(2 downto 0) := (others => '0');
   signal ldispCounter : unsigned(2 downto 0) := (others => '0');
   signal lastShift : std_logic := '0';
   signal lastState : std_logic := '0';
   signal state : unsigned(1 downto 0) := (others => '0');
   signal blank : std_logic := '0';

begin 
   process(clk50)
   begin
   --actually starts at counter = 1	  
      if rising_edge(clk50) then
         -- Count the lines and rows      
         if hCounter = hMaxCount-1 then
            hCounter <= (others => '0');
            if vCounter = vMaxCount-1 then
               vCounter <= (others => '0');
            else
               vCounter <= vCounter+1;
            end if;
         else
            hCounter <= hCounter+1;
         end if;

		 if hCounter = 39 or hCounter = 139 or hCounter = 239 or hCounter = 339 or hCounter = 439
		    or hCounter = 539 or hCounter = 639 or hCounter = 739 then
			hdispCounter <= hdispCounter + 1;
		 end if;
		 
		 if hCounter = 1 and (vCounter = 1 or vCounter = 75 or vCounter = 150 or vCounter = 225 or vCounter = 300
			or vCounter = 375 or vCounter = 450 or vCounter = 525) then
		    vdispCounter <= vdispCounter + 1;
		 end if;
		 
		 -- Are we in the display region?
		 if hCounter >= 40 and hCounter < 888 and vCounter >= 1 and vCounter < 601 then
			blank <= '0';
		 else 
			blank <= '1';
		 end if;
		 
         -- Are we in the hSync pulse?
         if hCounter >= hStartSync and hCounter < hEndSync then
            vga_hSync <= hsync_active;
         else
            vga_hSync <= not hsync_active;
         end if;

         -- Are we in the vSync pulse?
         if vCounter >= vStartSync and vCounter < vEndSync then
            vga_vSync <= vsync_active;
         else
            vga_vSync <= not vsync_active;
         end if;
		 
		 if blank = '0' then
			 if state = 0 then
				vga_red <= hdispCounter(0);
				vga_green <= hdispCounter(1);
				vga_blue <= hdispCounter(2);
			 elsif state = 1 then
				vga_red <= vdispCounter(0);
				vga_green <= vdispCounter(1);
				vga_blue <= vdispCounter(2);
			 else
				 if hCounter >= 239 and hCounter < 259 and vCounter >= 51 and vCounter < 251 then
					--I
					vga_red <= ldispCounter(0);
					vga_green <= ldispCounter(1);
					vga_blue <= ldispCounter(2);
				 elsif (vCounter = 51 and hCounter >= 583 and hCounter < 598) or (vCounter = 51 and hCounter >= 681 and hCounter < 696) or (vCounter = 52 and hCounter >= 580 and hCounter < 602) or (vCounter = 52 and hCounter >= 677 and hCounter < 699) or (vCounter = 53 and hCounter >= 577 and hCounter < 605) or (vCounter = 53 and hCounter >= 674 and hCounter < 702) or (vCounter = 54 and hCounter >= 576 and hCounter < 607) or (vCounter = 54 and hCounter >= 672 and hCounter < 703) or (vCounter = 55 and hCounter >= 574 and hCounter < 609) or (vCounter = 55 and hCounter >= 670 and hCounter < 705) or (vCounter = 56 and hCounter >= 573 and hCounter < 611) or (vCounter = 56 and hCounter >= 668 and hCounter < 706) or (vCounter = 57 and hCounter >= 572 and hCounter < 613) or (vCounter = 57 and hCounter >= 666 and hCounter < 707) or (vCounter = 58 and hCounter >= 571 and hCounter < 614) or (vCounter = 58 and hCounter >= 665 and hCounter < 708) or (vCounter = 59 and hCounter >= 570 and hCounter < 616) or (vCounter = 59 and hCounter >= 663 and hCounter < 709) or (vCounter = 60 and hCounter >= 569 and hCounter < 617) or (vCounter = 60 and hCounter >= 662 and hCounter < 710) or (vCounter = 61 and hCounter >= 568 and hCounter < 618) or (vCounter = 61 and hCounter >= 661 and hCounter < 711) or (vCounter = 62 and hCounter >= 567 and hCounter < 620) or (vCounter = 62 and hCounter >= 659 and hCounter < 712) or (vCounter = 63 and hCounter >= 567 and hCounter < 621) or (vCounter = 63 and hCounter >= 658 and hCounter < 712) or (vCounter = 64 and hCounter >= 566 and hCounter < 622) or (vCounter = 64 and hCounter >= 657 and hCounter < 713) or (vCounter = 65 and hCounter >= 565 and hCounter < 623) or (vCounter = 65 and hCounter >= 656 and hCounter < 714) or (vCounter = 66 and hCounter >= 565 and hCounter < 624) or (vCounter = 66 and hCounter >= 655 and hCounter < 714) or (vCounter = 67 and hCounter >= 564 and hCounter < 625) or (vCounter = 67 and hCounter >= 654 and hCounter < 715) or (vCounter = 68 and hCounter >= 564 and hCounter < 626) or (vCounter = 68 and hCounter >= 653 and hCounter < 715) or (vCounter = 69 and hCounter >= 563 and hCounter < 627) or (vCounter = 69 and hCounter >= 652 and hCounter < 716) or (vCounter = 70 and hCounter >= 563 and hCounter < 628) or (vCounter = 70 and hCounter >= 651 and hCounter < 716) or (vCounter = 71 and hCounter >= 563 and hCounter < 629) or (vCounter = 71 and hCounter >= 650 and hCounter < 716) or (vCounter = 72 and hCounter >= 562 and hCounter < 630) or (vCounter = 72 and hCounter >= 649 and hCounter < 717) or (vCounter = 73 and hCounter >= 562 and hCounter < 631) or (vCounter = 73 and hCounter >= 648 and hCounter < 717) or (vCounter = 74 and hCounter >= 562 and hCounter < 631) or (vCounter = 74 and hCounter >= 648 and hCounter < 717) or (vCounter = 75 and hCounter >= 561 and hCounter < 632) or (vCounter = 75 and hCounter >= 647 and hCounter < 718) or (vCounter = 76 and hCounter >= 561 and hCounter < 633) or (vCounter = 76 and hCounter >= 646 and hCounter < 718) or (vCounter = 77 and hCounter >= 561 and hCounter < 634) or (vCounter = 77 and hCounter >= 645 and hCounter < 718) or (vCounter = 78 and hCounter >= 561 and hCounter < 634) or (vCounter = 78 and hCounter >= 645 and hCounter < 718) or (vCounter = 79 and hCounter >= 561 and hCounter < 635) or (vCounter = 79 and hCounter >= 644 and hCounter < 718) or (vCounter = 80 and hCounter >= 560 and hCounter < 635) or (vCounter = 80 and hCounter >= 644 and hCounter < 719) or (vCounter = 81 and hCounter >= 560 and hCounter < 636) or (vCounter = 81 and hCounter >= 643 and hCounter < 719) or (vCounter = 82 and hCounter >= 560 and hCounter < 636) or (vCounter = 82 and hCounter >= 643 and hCounter < 719) or (vCounter = 83 and hCounter >= 560 and hCounter < 637) or (vCounter = 83 and hCounter >= 642 and hCounter < 719) or (vCounter = 84 and hCounter >= 560 and hCounter < 637) or (vCounter = 84 and hCounter >= 642 and hCounter < 719) or (vCounter = 85 and hCounter >= 560 and hCounter < 638) or (vCounter = 85 and hCounter >= 641 and hCounter < 719) or (vCounter = 86 and hCounter >= 560 and hCounter < 638) or (vCounter = 86 and hCounter >= 641 and hCounter < 719) or (vCounter = 87 and hCounter >= 560 and hCounter < 639) or (vCounter = 87 and hCounter >= 640 and hCounter < 719) or (vCounter = 88 and hCounter >= 560 and hCounter < 639) or (vCounter = 88 and hCounter >= 640 and hCounter < 719) or (vCounter = 89 and hCounter >= 560 and hCounter < 639) or (vCounter = 89 and hCounter >= 640 and hCounter < 719) or (vCounter = 90 and hCounter >= 560 and hCounter < 639) or (vCounter = 90 and hCounter >= 640 and hCounter < 719) or (vCounter = 91 and hCounter >= 560 and hCounter < 639) or (vCounter = 91 and hCounter >= 640 and hCounter < 719) or (vCounter = 92 and hCounter >= 560 and hCounter < 719) or (vCounter = 93 and hCounter >= 560 and hCounter < 719) or (vCounter = 94 and hCounter >= 560 and hCounter < 719) or (vCounter = 95 and hCounter >= 560 and hCounter < 719) or (vCounter = 96 and hCounter >= 560 and hCounter < 719) or (vCounter = 97 and hCounter >= 560 and hCounter < 719) or (vCounter = 98 and hCounter >= 560 and hCounter < 719) or (vCounter = 99 and hCounter >= 560 and hCounter < 719) or (vCounter = 100 and hCounter >= 560 and hCounter < 719) or (vCounter = 101 and hCounter >= 560 and hCounter < 719) or (vCounter = 102 and hCounter >= 560 and hCounter < 719) or (vCounter = 103 and hCounter >= 560 and hCounter < 719) or (vCounter = 104 and hCounter >= 560 and hCounter < 719) or (vCounter = 105 and hCounter >= 561 and hCounter < 718) or (vCounter = 106 and hCounter >= 561 and hCounter < 718) or (vCounter = 107 and hCounter >= 561 and hCounter < 718) or (vCounter = 108 and hCounter >= 561 and hCounter < 718) or (vCounter = 109 and hCounter >= 561 and hCounter < 718) or (vCounter = 110 and hCounter >= 561 and hCounter < 718) or (vCounter = 111 and hCounter >= 562 and hCounter < 717) or (vCounter = 112 and hCounter >= 562 and hCounter < 717) or (vCounter = 113 and hCounter >= 562 and hCounter < 717) or (vCounter = 114 and hCounter >= 562 and hCounter < 717) or (vCounter = 115 and hCounter >= 563 and hCounter < 716) or (vCounter = 116 and hCounter >= 563 and hCounter < 716) or (vCounter = 117 and hCounter >= 563 and hCounter < 716) or (vCounter = 118 and hCounter >= 563 and hCounter < 716) or (vCounter = 119 and hCounter >= 564 and hCounter < 715) or (vCounter = 120 and hCounter >= 564 and hCounter < 715) or (vCounter = 121 and hCounter >= 564 and hCounter < 715) or (vCounter = 122 and hCounter >= 564 and hCounter < 715) or (vCounter = 123 and hCounter >= 565 and hCounter < 714) or (vCounter = 124 and hCounter >= 565 and hCounter < 714) or (vCounter = 125 and hCounter >= 565 and hCounter < 714) or (vCounter = 126 and hCounter >= 566 and hCounter < 713) or (vCounter = 127 and hCounter >= 566 and hCounter < 713) or (vCounter = 128 and hCounter >= 566 and hCounter < 713) or (vCounter = 129 and hCounter >= 567 and hCounter < 712) or (vCounter = 130 and hCounter >= 567 and hCounter < 712) or (vCounter = 131 and hCounter >= 567 and hCounter < 712) or (vCounter = 132 and hCounter >= 568 and hCounter < 711) or (vCounter = 133 and hCounter >= 568 and hCounter < 711) or (vCounter = 134 and hCounter >= 569 and hCounter < 710) or (vCounter = 135 and hCounter >= 569 and hCounter < 710) or (vCounter = 136 and hCounter >= 569 and hCounter < 710) or (vCounter = 137 and hCounter >= 570 and hCounter < 709) or (vCounter = 138 and hCounter >= 570 and hCounter < 709) or (vCounter = 139 and hCounter >= 571 and hCounter < 708) or (vCounter = 140 and hCounter >= 571 and hCounter < 708) or (vCounter = 141 and hCounter >= 571 and hCounter < 708) or (vCounter = 142 and hCounter >= 572 and hCounter < 707) or (vCounter = 143 and hCounter >= 572 and hCounter < 707) or (vCounter = 144 and hCounter >= 573 and hCounter < 706) or (vCounter = 145 and hCounter >= 573 and hCounter < 706) or (vCounter = 146 and hCounter >= 574 and hCounter < 705) or (vCounter = 147 and hCounter >= 574 and hCounter < 705) or (vCounter = 148 and hCounter >= 575 and hCounter < 704) or (vCounter = 149 and hCounter >= 575 and hCounter < 704) or (vCounter = 150 and hCounter >= 575 and hCounter < 704) or (vCounter = 151 and hCounter >= 576 and hCounter < 703) or (vCounter = 152 and hCounter >= 576 and hCounter < 703) or (vCounter = 153 and hCounter >= 577 and hCounter < 702) or (vCounter = 154 and hCounter >= 577 and hCounter < 702) or (vCounter = 155 and hCounter >= 578 and hCounter < 701) or (vCounter = 156 and hCounter >= 579 and hCounter < 700) or (vCounter = 157 and hCounter >= 579 and hCounter < 700) or (vCounter = 158 and hCounter >= 580 and hCounter < 699) or (vCounter = 159 and hCounter >= 580 and hCounter < 699) or (vCounter = 160 and hCounter >= 581 and hCounter < 698) or (vCounter = 161 and hCounter >= 581 and hCounter < 698) or (vCounter = 162 and hCounter >= 582 and hCounter < 697) or (vCounter = 163 and hCounter >= 582 and hCounter < 697) or (vCounter = 164 and hCounter >= 583 and hCounter < 696) or (vCounter = 165 and hCounter >= 583 and hCounter < 696) or (vCounter = 166 and hCounter >= 584 and hCounter < 695) or (vCounter = 167 and hCounter >= 585 and hCounter < 694) or (vCounter = 168 and hCounter >= 585 and hCounter < 694) or (vCounter = 169 and hCounter >= 586 and hCounter < 693) or (vCounter = 170 and hCounter >= 586 and hCounter < 693) or (vCounter = 171 and hCounter >= 587 and hCounter < 692) or (vCounter = 172 and hCounter >= 588 and hCounter < 691) or (vCounter = 173 and hCounter >= 588 and hCounter < 691) or (vCounter = 174 and hCounter >= 589 and hCounter < 690) or (vCounter = 175 and hCounter >= 590 and hCounter < 689) or (vCounter = 176 and hCounter >= 590 and hCounter < 689) or (vCounter = 177 and hCounter >= 591 and hCounter < 688) or (vCounter = 178 and hCounter >= 591 and hCounter < 688) or (vCounter = 179 and hCounter >= 592 and hCounter < 687) or (vCounter = 180 and hCounter >= 593 and hCounter < 686) or (vCounter = 181 and hCounter >= 593 and hCounter < 686) or (vCounter = 182 and hCounter >= 594 and hCounter < 685) or (vCounter = 183 and hCounter >= 595 and hCounter < 684) or (vCounter = 184 and hCounter >= 595 and hCounter < 684) or (vCounter = 185 and hCounter >= 596 and hCounter < 683) or (vCounter = 186 and hCounter >= 597 and hCounter < 682) or (vCounter = 187 and hCounter >= 597 and hCounter < 682) or (vCounter = 188 and hCounter >= 598 and hCounter < 681) or (vCounter = 189 and hCounter >= 599 and hCounter < 680) or (vCounter = 190 and hCounter >= 600 and hCounter < 679) or (vCounter = 191 and hCounter >= 600 and hCounter < 679) or (vCounter = 192 and hCounter >= 601 and hCounter < 678) or (vCounter = 193 and hCounter >= 602 and hCounter < 677) or (vCounter = 194 and hCounter >= 602 and hCounter < 677) or (vCounter = 195 and hCounter >= 603 and hCounter < 676) or (vCounter = 196 and hCounter >= 604 and hCounter < 675) or (vCounter = 197 and hCounter >= 605 and hCounter < 674) or (vCounter = 198 and hCounter >= 605 and hCounter < 674) or (vCounter = 199 and hCounter >= 606 and hCounter < 673) or (vCounter = 200 and hCounter >= 607 and hCounter < 672) or (vCounter = 201 and hCounter >= 608 and hCounter < 671) or (vCounter = 202 and hCounter >= 608 and hCounter < 671) or (vCounter = 203 and hCounter >= 609 and hCounter < 670) or (vCounter = 204 and hCounter >= 610 and hCounter < 669) or (vCounter = 205 and hCounter >= 611 and hCounter < 668) or (vCounter = 206 and hCounter >= 611 and hCounter < 668) or (vCounter = 207 and hCounter >= 612 and hCounter < 667) or (vCounter = 208 and hCounter >= 613 and hCounter < 666) or (vCounter = 209 and hCounter >= 614 and hCounter < 665) or (vCounter = 210 and hCounter >= 614 and hCounter < 665) or (vCounter = 211 and hCounter >= 615 and hCounter < 664) or (vCounter = 212 and hCounter >= 616 and hCounter < 663) or (vCounter = 213 and hCounter >= 617 and hCounter < 662) or (vCounter = 214 and hCounter >= 617 and hCounter < 662) or (vCounter = 215 and hCounter >= 618 and hCounter < 661) or (vCounter = 216 and hCounter >= 619 and hCounter < 660) or (vCounter = 217 and hCounter >= 620 and hCounter < 659) or (vCounter = 218 and hCounter >= 620 and hCounter < 659) or (vCounter = 219 and hCounter >= 621 and hCounter < 658) or (vCounter = 220 and hCounter >= 622 and hCounter < 657) or (vCounter = 221 and hCounter >= 623 and hCounter < 656) or (vCounter = 222 and hCounter >= 623 and hCounter < 656) or (vCounter = 223 and hCounter >= 624 and hCounter < 655) or (vCounter = 224 and hCounter >= 625 and hCounter < 654) or (vCounter = 225 and hCounter >= 626 and hCounter < 653) or (vCounter = 226 and hCounter >= 626 and hCounter < 653) or (vCounter = 227 and hCounter >= 627 and hCounter < 652) or (vCounter = 228 and hCounter >= 628 and hCounter < 651) or (vCounter = 229 and hCounter >= 629 and hCounter < 650) or (vCounter = 230 and hCounter >= 629 and hCounter < 650) or (vCounter = 231 and hCounter >= 630 and hCounter < 649) or (vCounter = 232 and hCounter >= 631 and hCounter < 648) or (vCounter = 233 and hCounter >= 631 and hCounter < 648) or (vCounter = 234 and hCounter >= 632 and hCounter < 647) or (vCounter = 235 and hCounter >= 633 and hCounter < 646) or (vCounter = 236 and hCounter >= 633 and hCounter < 646) or (vCounter = 237 and hCounter >= 634 and hCounter < 645) or (vCounter = 238 and hCounter >= 634 and hCounter < 645) or (vCounter = 239 and hCounter >= 635 and hCounter < 644) or (vCounter = 240 and hCounter >= 635 and hCounter < 644) or (vCounter = 241 and hCounter >= 636 and hCounter < 643) or (vCounter = 242 and hCounter >= 637 and hCounter < 642) or (vCounter = 243 and hCounter >= 637 and hCounter < 642) or (vCounter = 244 and hCounter >= 637 and hCounter < 642) or (vCounter = 245 and hCounter >= 638 and hCounter < 641) or (vCounter = 246 and hCounter >= 638 and hCounter < 641) or (vCounter = 247 and hCounter >= 639 and hCounter < 640) or (vCounter = 248 and hCounter >= 639 and hCounter < 640) or (vCounter = 249 and hCounter >= 639 and hCounter < 640) or (vCounter = 250 and hCounter >= 639 and hCounter < 640) then
					--?
					vga_red <= ldispCounter(0);
					vga_green <= ldispCounter(1);
					vga_blue <= ldispCounter(2);
				 elsif (vCounter = 351 and hCounter >= 140 and hCounter < 159) or (vCounter = 351 and hCounter >= 220 and hCounter < 239) or (vCounter = 352 and hCounter >= 140 and hCounter < 160) or (vCounter = 352 and hCounter >= 219 and hCounter < 239) or (vCounter = 353 and hCounter >= 140 and hCounter < 160) or (vCounter = 353 and hCounter >= 219 and hCounter < 239) or (vCounter = 354 and hCounter >= 140 and hCounter < 160) or (vCounter = 354 and hCounter >= 219 and hCounter < 239) or (vCounter = 355 and hCounter >= 140 and hCounter < 160) or (vCounter = 355 and hCounter >= 219 and hCounter < 239) or (vCounter = 356 and hCounter >= 141 and hCounter < 160) or (vCounter = 356 and hCounter >= 219 and hCounter < 238) or (vCounter = 357 and hCounter >= 141 and hCounter < 161) or (vCounter = 357 and hCounter >= 218 and hCounter < 238) or (vCounter = 358 and hCounter >= 141 and hCounter < 161) or (vCounter = 358 and hCounter >= 218 and hCounter < 238) or (vCounter = 359 and hCounter >= 141 and hCounter < 161) or (vCounter = 359 and hCounter >= 218 and hCounter < 238) or (vCounter = 360 and hCounter >= 141 and hCounter < 161) or (vCounter = 360 and hCounter >= 218 and hCounter < 238) or (vCounter = 361 and hCounter >= 142 and hCounter < 161) or (vCounter = 361 and hCounter >= 218 and hCounter < 237) or (vCounter = 362 and hCounter >= 142 and hCounter < 162) or (vCounter = 362 and hCounter >= 217 and hCounter < 237) or (vCounter = 363 and hCounter >= 142 and hCounter < 162) or (vCounter = 363 and hCounter >= 217 and hCounter < 237) or (vCounter = 364 and hCounter >= 142 and hCounter < 162) or (vCounter = 364 and hCounter >= 217 and hCounter < 237) or (vCounter = 365 and hCounter >= 142 and hCounter < 162) or (vCounter = 365 and hCounter >= 217 and hCounter < 237) or (vCounter = 366 and hCounter >= 143 and hCounter < 162) or (vCounter = 366 and hCounter >= 217 and hCounter < 236) or (vCounter = 367 and hCounter >= 143 and hCounter < 163) or (vCounter = 367 and hCounter >= 216 and hCounter < 236) or (vCounter = 368 and hCounter >= 143 and hCounter < 163) or (vCounter = 368 and hCounter >= 216 and hCounter < 236) or (vCounter = 369 and hCounter >= 143 and hCounter < 163) or (vCounter = 369 and hCounter >= 216 and hCounter < 236) or (vCounter = 370 and hCounter >= 143 and hCounter < 163) or (vCounter = 370 and hCounter >= 216 and hCounter < 236) or (vCounter = 371 and hCounter >= 144 and hCounter < 163) or (vCounter = 371 and hCounter >= 216 and hCounter < 235) or (vCounter = 372 and hCounter >= 144 and hCounter < 164) or (vCounter = 372 and hCounter >= 215 and hCounter < 235) or (vCounter = 373 and hCounter >= 144 and hCounter < 164) or (vCounter = 373 and hCounter >= 215 and hCounter < 235) or (vCounter = 374 and hCounter >= 144 and hCounter < 164) or (vCounter = 374 and hCounter >= 215 and hCounter < 235) or (vCounter = 375 and hCounter >= 144 and hCounter < 164) or (vCounter = 375 and hCounter >= 215 and hCounter < 235) or (vCounter = 376 and hCounter >= 145 and hCounter < 164) or (vCounter = 376 and hCounter >= 215 and hCounter < 234) or (vCounter = 377 and hCounter >= 145 and hCounter < 165) or (vCounter = 377 and hCounter >= 214 and hCounter < 234) or (vCounter = 378 and hCounter >= 145 and hCounter < 165) or (vCounter = 378 and hCounter >= 214 and hCounter < 234) or (vCounter = 379 and hCounter >= 145 and hCounter < 165) or (vCounter = 379 and hCounter >= 214 and hCounter < 234) or (vCounter = 380 and hCounter >= 145 and hCounter < 165) or (vCounter = 380 and hCounter >= 214 and hCounter < 234) or (vCounter = 381 and hCounter >= 146 and hCounter < 165) or (vCounter = 381 and hCounter >= 214 and hCounter < 233) or (vCounter = 382 and hCounter >= 146 and hCounter < 166) or (vCounter = 382 and hCounter >= 213 and hCounter < 233) or (vCounter = 383 and hCounter >= 146 and hCounter < 166) or (vCounter = 383 and hCounter >= 213 and hCounter < 233) or (vCounter = 384 and hCounter >= 146 and hCounter < 166) or (vCounter = 384 and hCounter >= 213 and hCounter < 233) or (vCounter = 385 and hCounter >= 146 and hCounter < 166) or (vCounter = 385 and hCounter >= 213 and hCounter < 233) or (vCounter = 386 and hCounter >= 147 and hCounter < 166) or (vCounter = 386 and hCounter >= 213 and hCounter < 232) or (vCounter = 387 and hCounter >= 147 and hCounter < 167) or (vCounter = 387 and hCounter >= 212 and hCounter < 232) or (vCounter = 388 and hCounter >= 147 and hCounter < 167) or (vCounter = 388 and hCounter >= 212 and hCounter < 232) or (vCounter = 389 and hCounter >= 147 and hCounter < 167) or (vCounter = 389 and hCounter >= 212 and hCounter < 232) or (vCounter = 390 and hCounter >= 147 and hCounter < 167) or (vCounter = 390 and hCounter >= 212 and hCounter < 232) or (vCounter = 391 and hCounter >= 148 and hCounter < 167) or (vCounter = 391 and hCounter >= 212 and hCounter < 231) or (vCounter = 392 and hCounter >= 148 and hCounter < 168) or (vCounter = 392 and hCounter >= 211 and hCounter < 231) or (vCounter = 393 and hCounter >= 148 and hCounter < 168) or (vCounter = 393 and hCounter >= 211 and hCounter < 231) or (vCounter = 394 and hCounter >= 148 and hCounter < 168) or (vCounter = 394 and hCounter >= 211 and hCounter < 231) or (vCounter = 395 and hCounter >= 148 and hCounter < 168) or (vCounter = 395 and hCounter >= 211 and hCounter < 231) or (vCounter = 396 and hCounter >= 149 and hCounter < 168) or (vCounter = 396 and hCounter >= 211 and hCounter < 230) or (vCounter = 397 and hCounter >= 149 and hCounter < 169) or (vCounter = 397 and hCounter >= 210 and hCounter < 230) or (vCounter = 398 and hCounter >= 149 and hCounter < 169) or (vCounter = 398 and hCounter >= 210 and hCounter < 230) or (vCounter = 399 and hCounter >= 149 and hCounter < 169) or (vCounter = 399 and hCounter >= 210 and hCounter < 230) or (vCounter = 400 and hCounter >= 149 and hCounter < 169) or (vCounter = 400 and hCounter >= 210 and hCounter < 230) or (vCounter = 401 and hCounter >= 150 and hCounter < 169) or (vCounter = 401 and hCounter >= 210 and hCounter < 229) or (vCounter = 402 and hCounter >= 150 and hCounter < 170) or (vCounter = 402 and hCounter >= 209 and hCounter < 229) or (vCounter = 403 and hCounter >= 150 and hCounter < 170) or (vCounter = 403 and hCounter >= 209 and hCounter < 229) or (vCounter = 404 and hCounter >= 150 and hCounter < 170) or (vCounter = 404 and hCounter >= 209 and hCounter < 229) or (vCounter = 405 and hCounter >= 150 and hCounter < 170) or (vCounter = 405 and hCounter >= 209 and hCounter < 229) or (vCounter = 406 and hCounter >= 151 and hCounter < 170) or (vCounter = 406 and hCounter >= 209 and hCounter < 228) or (vCounter = 407 and hCounter >= 151 and hCounter < 171) or (vCounter = 407 and hCounter >= 208 and hCounter < 228) or (vCounter = 408 and hCounter >= 151 and hCounter < 171) or (vCounter = 408 and hCounter >= 208 and hCounter < 228) or (vCounter = 409 and hCounter >= 151 and hCounter < 171) or (vCounter = 409 and hCounter >= 208 and hCounter < 228) or (vCounter = 410 and hCounter >= 151 and hCounter < 171) or (vCounter = 410 and hCounter >= 208 and hCounter < 228) or (vCounter = 411 and hCounter >= 152 and hCounter < 171) or (vCounter = 411 and hCounter >= 208 and hCounter < 227) or (vCounter = 412 and hCounter >= 152 and hCounter < 172) or (vCounter = 412 and hCounter >= 207 and hCounter < 227) or (vCounter = 413 and hCounter >= 152 and hCounter < 172) or (vCounter = 413 and hCounter >= 207 and hCounter < 227) or (vCounter = 414 and hCounter >= 152 and hCounter < 172) or (vCounter = 414 and hCounter >= 207 and hCounter < 227) or (vCounter = 415 and hCounter >= 152 and hCounter < 172) or (vCounter = 415 and hCounter >= 207 and hCounter < 227) or (vCounter = 416 and hCounter >= 153 and hCounter < 172) or (vCounter = 416 and hCounter >= 207 and hCounter < 226) or (vCounter = 417 and hCounter >= 153 and hCounter < 173) or (vCounter = 417 and hCounter >= 206 and hCounter < 226) or (vCounter = 418 and hCounter >= 153 and hCounter < 173) or (vCounter = 418 and hCounter >= 206 and hCounter < 226) or (vCounter = 419 and hCounter >= 153 and hCounter < 173) or (vCounter = 419 and hCounter >= 206 and hCounter < 226) or (vCounter = 420 and hCounter >= 153 and hCounter < 173) or (vCounter = 420 and hCounter >= 206 and hCounter < 226) or (vCounter = 421 and hCounter >= 154 and hCounter < 173) or (vCounter = 421 and hCounter >= 206 and hCounter < 225) or (vCounter = 422 and hCounter >= 154 and hCounter < 174) or (vCounter = 422 and hCounter >= 205 and hCounter < 225) or (vCounter = 423 and hCounter >= 154 and hCounter < 174) or (vCounter = 423 and hCounter >= 205 and hCounter < 225) or (vCounter = 424 and hCounter >= 154 and hCounter < 174) or (vCounter = 424 and hCounter >= 205 and hCounter < 225) or (vCounter = 425 and hCounter >= 154 and hCounter < 174) or (vCounter = 425 and hCounter >= 205 and hCounter < 225) or (vCounter = 426 and hCounter >= 155 and hCounter < 174) or (vCounter = 426 and hCounter >= 205 and hCounter < 224) or (vCounter = 427 and hCounter >= 155 and hCounter < 175) or (vCounter = 427 and hCounter >= 204 and hCounter < 224) or (vCounter = 428 and hCounter >= 155 and hCounter < 175) or (vCounter = 428 and hCounter >= 204 and hCounter < 224) or (vCounter = 429 and hCounter >= 155 and hCounter < 175) or (vCounter = 429 and hCounter >= 204 and hCounter < 224) or (vCounter = 430 and hCounter >= 155 and hCounter < 175) or (vCounter = 430 and hCounter >= 204 and hCounter < 224) or (vCounter = 431 and hCounter >= 156 and hCounter < 175) or (vCounter = 431 and hCounter >= 204 and hCounter < 223) or (vCounter = 432 and hCounter >= 156 and hCounter < 176) or (vCounter = 432 and hCounter >= 203 and hCounter < 223) or (vCounter = 433 and hCounter >= 156 and hCounter < 176) or (vCounter = 433 and hCounter >= 203 and hCounter < 223) or (vCounter = 434 and hCounter >= 156 and hCounter < 176) or (vCounter = 434 and hCounter >= 203 and hCounter < 223) or (vCounter = 435 and hCounter >= 156 and hCounter < 176) or (vCounter = 435 and hCounter >= 203 and hCounter < 223) or (vCounter = 436 and hCounter >= 157 and hCounter < 176) or (vCounter = 436 and hCounter >= 203 and hCounter < 222) or (vCounter = 437 and hCounter >= 157 and hCounter < 177) or (vCounter = 437 and hCounter >= 202 and hCounter < 222) or (vCounter = 438 and hCounter >= 157 and hCounter < 177) or (vCounter = 438 and hCounter >= 202 and hCounter < 222) or (vCounter = 439 and hCounter >= 157 and hCounter < 177) or (vCounter = 439 and hCounter >= 202 and hCounter < 222) or (vCounter = 440 and hCounter >= 157 and hCounter < 177) or (vCounter = 440 and hCounter >= 202 and hCounter < 222) or (vCounter = 441 and hCounter >= 158 and hCounter < 177) or (vCounter = 441 and hCounter >= 202 and hCounter < 221) or (vCounter = 442 and hCounter >= 158 and hCounter < 178) or (vCounter = 442 and hCounter >= 201 and hCounter < 221) or (vCounter = 443 and hCounter >= 158 and hCounter < 178) or (vCounter = 443 and hCounter >= 201 and hCounter < 221) or (vCounter = 444 and hCounter >= 158 and hCounter < 178) or (vCounter = 444 and hCounter >= 201 and hCounter < 221) or (vCounter = 445 and hCounter >= 158 and hCounter < 178) or (vCounter = 445 and hCounter >= 201 and hCounter < 221) or (vCounter = 446 and hCounter >= 159 and hCounter < 178) or (vCounter = 446 and hCounter >= 201 and hCounter < 220) or (vCounter = 447 and hCounter >= 159 and hCounter < 179) or (vCounter = 447 and hCounter >= 200 and hCounter < 220) or (vCounter = 448 and hCounter >= 159 and hCounter < 179) or (vCounter = 448 and hCounter >= 200 and hCounter < 220) or (vCounter = 449 and hCounter >= 159 and hCounter < 179) or (vCounter = 449 and hCounter >= 200 and hCounter < 220) or (vCounter = 450 and hCounter >= 159 and hCounter < 179) or (vCounter = 450 and hCounter >= 200 and hCounter < 220) or (vCounter = 451 and hCounter >= 160 and hCounter < 179) or (vCounter = 451 and hCounter >= 200 and hCounter < 219) or (vCounter = 452 and hCounter >= 160 and hCounter < 180) or (vCounter = 452 and hCounter >= 199 and hCounter < 219) or (vCounter = 453 and hCounter >= 160 and hCounter < 180) or (vCounter = 453 and hCounter >= 199 and hCounter < 219) or (vCounter = 454 and hCounter >= 160 and hCounter < 180) or (vCounter = 454 and hCounter >= 199 and hCounter < 219) or (vCounter = 455 and hCounter >= 160 and hCounter < 180) or (vCounter = 455 and hCounter >= 199 and hCounter < 219) or (vCounter = 456 and hCounter >= 161 and hCounter < 180) or (vCounter = 456 and hCounter >= 199 and hCounter < 218) or (vCounter = 457 and hCounter >= 161 and hCounter < 181) or (vCounter = 457 and hCounter >= 198 and hCounter < 218) or (vCounter = 458 and hCounter >= 161 and hCounter < 181) or (vCounter = 458 and hCounter >= 198 and hCounter < 218) or (vCounter = 459 and hCounter >= 161 and hCounter < 181) or (vCounter = 459 and hCounter >= 198 and hCounter < 218) or (vCounter = 460 and hCounter >= 161 and hCounter < 181) or (vCounter = 460 and hCounter >= 198 and hCounter < 218) or (vCounter = 461 and hCounter >= 162 and hCounter < 181) or (vCounter = 461 and hCounter >= 198 and hCounter < 217) or (vCounter = 462 and hCounter >= 162 and hCounter < 182) or (vCounter = 462 and hCounter >= 197 and hCounter < 217) or (vCounter = 463 and hCounter >= 162 and hCounter < 182) or (vCounter = 463 and hCounter >= 197 and hCounter < 217) or (vCounter = 464 and hCounter >= 162 and hCounter < 182) or (vCounter = 464 and hCounter >= 197 and hCounter < 217) or (vCounter = 465 and hCounter >= 162 and hCounter < 182) or (vCounter = 465 and hCounter >= 197 and hCounter < 217) or (vCounter = 466 and hCounter >= 163 and hCounter < 182) or (vCounter = 466 and hCounter >= 197 and hCounter < 216) or (vCounter = 467 and hCounter >= 163 and hCounter < 183) or (vCounter = 467 and hCounter >= 196 and hCounter < 216) or (vCounter = 468 and hCounter >= 163 and hCounter < 183) or (vCounter = 468 and hCounter >= 196 and hCounter < 216) or (vCounter = 469 and hCounter >= 163 and hCounter < 183) or (vCounter = 469 and hCounter >= 196 and hCounter < 216) or (vCounter = 470 and hCounter >= 163 and hCounter < 183) or (vCounter = 470 and hCounter >= 196 and hCounter < 216) or (vCounter = 471 and hCounter >= 164 and hCounter < 183) or (vCounter = 471 and hCounter >= 196 and hCounter < 215) or (vCounter = 472 and hCounter >= 164 and hCounter < 184) or (vCounter = 472 and hCounter >= 195 and hCounter < 215) or (vCounter = 473 and hCounter >= 164 and hCounter < 184) or (vCounter = 473 and hCounter >= 195 and hCounter < 215) or (vCounter = 474 and hCounter >= 164 and hCounter < 184) or (vCounter = 474 and hCounter >= 195 and hCounter < 215) or (vCounter = 475 and hCounter >= 164 and hCounter < 184) or (vCounter = 475 and hCounter >= 195 and hCounter < 215) or (vCounter = 476 and hCounter >= 165 and hCounter < 184) or (vCounter = 476 and hCounter >= 195 and hCounter < 214) or (vCounter = 477 and hCounter >= 165 and hCounter < 185) or (vCounter = 477 and hCounter >= 194 and hCounter < 214) or (vCounter = 478 and hCounter >= 165 and hCounter < 185) or (vCounter = 478 and hCounter >= 194 and hCounter < 214) or (vCounter = 479 and hCounter >= 165 and hCounter < 185) or (vCounter = 479 and hCounter >= 194 and hCounter < 214) or (vCounter = 480 and hCounter >= 165 and hCounter < 185) or (vCounter = 480 and hCounter >= 194 and hCounter < 214) or (vCounter = 481 and hCounter >= 166 and hCounter < 185) or (vCounter = 481 and hCounter >= 194 and hCounter < 213) or (vCounter = 482 and hCounter >= 166 and hCounter < 186) or (vCounter = 482 and hCounter >= 193 and hCounter < 213) or (vCounter = 483 and hCounter >= 166 and hCounter < 186) or (vCounter = 483 and hCounter >= 193 and hCounter < 213) or (vCounter = 484 and hCounter >= 166 and hCounter < 186) or (vCounter = 484 and hCounter >= 193 and hCounter < 213) or (vCounter = 485 and hCounter >= 166 and hCounter < 186) or (vCounter = 485 and hCounter >= 193 and hCounter < 213) or (vCounter = 486 and hCounter >= 167 and hCounter < 186) or (vCounter = 486 and hCounter >= 193 and hCounter < 212) or (vCounter = 487 and hCounter >= 167 and hCounter < 187) or (vCounter = 487 and hCounter >= 192 and hCounter < 212) or (vCounter = 488 and hCounter >= 167 and hCounter < 187) or (vCounter = 488 and hCounter >= 192 and hCounter < 212) or (vCounter = 489 and hCounter >= 167 and hCounter < 187) or (vCounter = 489 and hCounter >= 192 and hCounter < 212) or (vCounter = 490 and hCounter >= 167 and hCounter < 187) or (vCounter = 490 and hCounter >= 192 and hCounter < 212) or (vCounter = 491 and hCounter >= 168 and hCounter < 187) or (vCounter = 491 and hCounter >= 192 and hCounter < 211) or (vCounter = 492 and hCounter >= 168 and hCounter < 188) or (vCounter = 492 and hCounter >= 191 and hCounter < 211) or (vCounter = 493 and hCounter >= 168 and hCounter < 188) or (vCounter = 493 and hCounter >= 191 and hCounter < 211) or (vCounter = 494 and hCounter >= 168 and hCounter < 188) or (vCounter = 494 and hCounter >= 191 and hCounter < 211) or (vCounter = 495 and hCounter >= 168 and hCounter < 188) or (vCounter = 495 and hCounter >= 191 and hCounter < 211) or (vCounter = 496 and hCounter >= 169 and hCounter < 188) or (vCounter = 496 and hCounter >= 191 and hCounter < 210) or (vCounter = 497 and hCounter >= 169 and hCounter < 189) or (vCounter = 497 and hCounter >= 190 and hCounter < 210) or (vCounter = 498 and hCounter >= 169 and hCounter < 189) or (vCounter = 498 and hCounter >= 190 and hCounter < 210) or (vCounter = 499 and hCounter >= 169 and hCounter < 189) or (vCounter = 499 and hCounter >= 190 and hCounter < 210) or (vCounter = 500 and hCounter >= 169 and hCounter < 189) or (vCounter = 500 and hCounter >= 190 and hCounter < 210) or (vCounter = 501 and hCounter >= 170 and hCounter < 189) or (vCounter = 501 and hCounter >= 190 and hCounter < 209) or (vCounter = 502 and hCounter >= 170 and hCounter < 209) or (vCounter = 503 and hCounter >= 170 and hCounter < 209) or (vCounter = 504 and hCounter >= 170 and hCounter < 209) or (vCounter = 505 and hCounter >= 170 and hCounter < 209) or (vCounter = 506 and hCounter >= 171 and hCounter < 208) or (vCounter = 507 and hCounter >= 171 and hCounter < 208) or (vCounter = 508 and hCounter >= 171 and hCounter < 208) or (vCounter = 509 and hCounter >= 171 and hCounter < 208) or (vCounter = 510 and hCounter >= 171 and hCounter < 208) or (vCounter = 511 and hCounter >= 172 and hCounter < 207) or (vCounter = 512 and hCounter >= 172 and hCounter < 207) or (vCounter = 513 and hCounter >= 172 and hCounter < 207) or (vCounter = 514 and hCounter >= 172 and hCounter < 207) or (vCounter = 515 and hCounter >= 172 and hCounter < 207) or (vCounter = 516 and hCounter >= 173 and hCounter < 206) or (vCounter = 517 and hCounter >= 173 and hCounter < 206) or (vCounter = 518 and hCounter >= 173 and hCounter < 206) or (vCounter = 519 and hCounter >= 173 and hCounter < 206) or (vCounter = 520 and hCounter >= 173 and hCounter < 206) or (vCounter = 521 and hCounter >= 174 and hCounter < 205) or (vCounter = 522 and hCounter >= 174 and hCounter < 205) or (vCounter = 523 and hCounter >= 174 and hCounter < 205) or (vCounter = 524 and hCounter >= 174 and hCounter < 205) or (vCounter = 525 and hCounter >= 174 and hCounter < 205) or (vCounter = 526 and hCounter >= 175 and hCounter < 204) or (vCounter = 527 and hCounter >= 175 and hCounter < 204) or (vCounter = 528 and hCounter >= 175 and hCounter < 204) or (vCounter = 529 and hCounter >= 175 and hCounter < 204) or (vCounter = 530 and hCounter >= 175 and hCounter < 204) or (vCounter = 531 and hCounter >= 176 and hCounter < 203) or (vCounter = 532 and hCounter >= 176 and hCounter < 203) or (vCounter = 533 and hCounter >= 176 and hCounter < 203) or (vCounter = 534 and hCounter >= 176 and hCounter < 203) or (vCounter = 535 and hCounter >= 176 and hCounter < 203) or (vCounter = 536 and hCounter >= 177 and hCounter < 202) or (vCounter = 537 and hCounter >= 177 and hCounter < 202) or (vCounter = 538 and hCounter >= 177 and hCounter < 202) or (vCounter = 539 and hCounter >= 177 and hCounter < 202) or (vCounter = 540 and hCounter >= 177 and hCounter < 202) or (vCounter = 541 and hCounter >= 178 and hCounter < 201) or (vCounter = 542 and hCounter >= 178 and hCounter < 201) or (vCounter = 543 and hCounter >= 178 and hCounter < 201) or (vCounter = 544 and hCounter >= 178 and hCounter < 201) or (vCounter = 545 and hCounter >= 178 and hCounter < 201) or (vCounter = 546 and hCounter >= 179 and hCounter < 200) or (vCounter = 547 and hCounter >= 179 and hCounter < 200) or (vCounter = 548 and hCounter >= 179 and hCounter < 200) or (vCounter = 549 and hCounter >= 179 and hCounter < 200) or (vCounter = 550 and hCounter >= 179 and hCounter < 200) then
					--V
					vga_red <= ldispCounter(0);
					vga_green <= ldispCounter(1);
					vga_blue <= ldispCounter(2);
				 elsif (hCounter > 339 and hCounter <= 359 and vCounter > 351 and vCounter < 551) or (hCounter > 419 and hCounter <= 439 and vCounter > 351 and vCounter < 551) or (hCounter > 339 and hCounter < 439 and vCounter > 441 and vCounter < 461) then
					--H
					vga_red <= ldispCounter(0);
					vga_green <= ldispCounter(1);
					vga_blue <= ldispCounter(2);
				 elsif (vCounter = 351 and hCounter >= 520 and hCounter < 539) or (vCounter = 352 and hCounter >= 520 and hCounter < 554) or (vCounter = 353 and hCounter >= 520 and hCounter < 559) or (vCounter = 354 and hCounter >= 520 and hCounter < 564) or (vCounter = 355 and hCounter >= 520 and hCounter < 567) or (vCounter = 356 and hCounter >= 520 and hCounter < 571) or (vCounter = 357 and hCounter >= 520 and hCounter < 574) or (vCounter = 358 and hCounter >= 520 and hCounter < 576) or (vCounter = 359 and hCounter >= 520 and hCounter < 579) or (vCounter = 360 and hCounter >= 520 and hCounter < 581) or (vCounter = 361 and hCounter >= 520 and hCounter < 583) or (vCounter = 362 and hCounter >= 520 and hCounter < 585) or (vCounter = 363 and hCounter >= 520 and hCounter < 587) or (vCounter = 364 and hCounter >= 520 and hCounter < 589) or (vCounter = 365 and hCounter >= 520 and hCounter < 591) or (vCounter = 366 and hCounter >= 520 and hCounter < 592) or (vCounter = 367 and hCounter >= 520 and hCounter < 594) or (vCounter = 368 and hCounter >= 520 and hCounter < 595) or (vCounter = 369 and hCounter >= 520 and hCounter < 597) or (vCounter = 370 and hCounter >= 520 and hCounter < 598) or (vCounter = 371 and hCounter >= 520 and hCounter < 539) or (vCounter = 371 and hCounter >= 540 and hCounter < 599) or (vCounter = 372 and hCounter >= 520 and hCounter < 539) or (vCounter = 372 and hCounter >= 552 and hCounter < 601) or (vCounter = 373 and hCounter >= 520 and hCounter < 539) or (vCounter = 373 and hCounter >= 557 and hCounter < 602) or (vCounter = 374 and hCounter >= 520 and hCounter < 539) or (vCounter = 374 and hCounter >= 561 and hCounter < 603) or (vCounter = 375 and hCounter >= 520 and hCounter < 539) or (vCounter = 375 and hCounter >= 564 and hCounter < 604) or (vCounter = 376 and hCounter >= 520 and hCounter < 539) or (vCounter = 376 and hCounter >= 567 and hCounter < 606) or (vCounter = 377 and hCounter >= 520 and hCounter < 539) or (vCounter = 377 and hCounter >= 570 and hCounter < 607) or (vCounter = 378 and hCounter >= 520 and hCounter < 539) or (vCounter = 378 and hCounter >= 572 and hCounter < 608) or (vCounter = 379 and hCounter >= 520 and hCounter < 539) or (vCounter = 379 and hCounter >= 574 and hCounter < 609) or (vCounter = 380 and hCounter >= 520 and hCounter < 539) or (vCounter = 380 and hCounter >= 576 and hCounter < 610) or (vCounter = 381 and hCounter >= 520 and hCounter < 539) or (vCounter = 381 and hCounter >= 578 and hCounter < 611) or (vCounter = 382 and hCounter >= 520 and hCounter < 539) or (vCounter = 382 and hCounter >= 580 and hCounter < 612) or (vCounter = 383 and hCounter >= 520 and hCounter < 539) or (vCounter = 383 and hCounter >= 582 and hCounter < 613) or (vCounter = 384 and hCounter >= 520 and hCounter < 539) or (vCounter = 384 and hCounter >= 583 and hCounter < 614) or (vCounter = 385 and hCounter >= 520 and hCounter < 539) or (vCounter = 385 and hCounter >= 585 and hCounter < 615) or (vCounter = 386 and hCounter >= 520 and hCounter < 539) or (vCounter = 386 and hCounter >= 586 and hCounter < 615) or (vCounter = 387 and hCounter >= 520 and hCounter < 539) or (vCounter = 387 and hCounter >= 588 and hCounter < 616) or (vCounter = 388 and hCounter >= 520 and hCounter < 539) or (vCounter = 388 and hCounter >= 589 and hCounter < 617) or (vCounter = 389 and hCounter >= 520 and hCounter < 539) or (vCounter = 389 and hCounter >= 590 and hCounter < 618) or (vCounter = 390 and hCounter >= 520 and hCounter < 539) or (vCounter = 390 and hCounter >= 591 and hCounter < 619) or (vCounter = 391 and hCounter >= 520 and hCounter < 539) or (vCounter = 391 and hCounter >= 592 and hCounter < 619) or (vCounter = 392 and hCounter >= 520 and hCounter < 539) or (vCounter = 392 and hCounter >= 594 and hCounter < 620) or (vCounter = 393 and hCounter >= 520 and hCounter < 539) or (vCounter = 393 and hCounter >= 595 and hCounter < 621) or (vCounter = 394 and hCounter >= 520 and hCounter < 539) or (vCounter = 394 and hCounter >= 596 and hCounter < 622) or (vCounter = 395 and hCounter >= 520 and hCounter < 539) or (vCounter = 395 and hCounter >= 597 and hCounter < 622) or (vCounter = 396 and hCounter >= 520 and hCounter < 539) or (vCounter = 396 and hCounter >= 598 and hCounter < 623) or (vCounter = 397 and hCounter >= 520 and hCounter < 539) or (vCounter = 397 and hCounter >= 599 and hCounter < 624) or (vCounter = 398 and hCounter >= 520 and hCounter < 539) or (vCounter = 398 and hCounter >= 599 and hCounter < 624) or (vCounter = 399 and hCounter >= 520 and hCounter < 539) or (vCounter = 399 and hCounter >= 600 and hCounter < 625) or (vCounter = 400 and hCounter >= 520 and hCounter < 539) or (vCounter = 400 and hCounter >= 601 and hCounter < 626) or (vCounter = 401 and hCounter >= 520 and hCounter < 539) or (vCounter = 401 and hCounter >= 602 and hCounter < 626) or (vCounter = 402 and hCounter >= 520 and hCounter < 539) or (vCounter = 402 and hCounter >= 603 and hCounter < 627) or (vCounter = 403 and hCounter >= 520 and hCounter < 539) or (vCounter = 403 and hCounter >= 604 and hCounter < 627) or (vCounter = 404 and hCounter >= 520 and hCounter < 539) or (vCounter = 404 and hCounter >= 604 and hCounter < 628) or (vCounter = 405 and hCounter >= 520 and hCounter < 539) or (vCounter = 405 and hCounter >= 605 and hCounter < 628) or (vCounter = 406 and hCounter >= 520 and hCounter < 539) or (vCounter = 406 and hCounter >= 606 and hCounter < 629) or (vCounter = 407 and hCounter >= 520 and hCounter < 539) or (vCounter = 407 and hCounter >= 606 and hCounter < 629) or (vCounter = 408 and hCounter >= 520 and hCounter < 539) or (vCounter = 408 and hCounter >= 607 and hCounter < 630) or (vCounter = 409 and hCounter >= 520 and hCounter < 539) or (vCounter = 409 and hCounter >= 608 and hCounter < 630) or (vCounter = 410 and hCounter >= 520 and hCounter < 539) or (vCounter = 410 and hCounter >= 608 and hCounter < 631) or (vCounter = 411 and hCounter >= 520 and hCounter < 539) or (vCounter = 411 and hCounter >= 609 and hCounter < 631) or (vCounter = 412 and hCounter >= 520 and hCounter < 539) or (vCounter = 412 and hCounter >= 609 and hCounter < 632) or (vCounter = 413 and hCounter >= 520 and hCounter < 539) or (vCounter = 413 and hCounter >= 610 and hCounter < 632) or (vCounter = 414 and hCounter >= 520 and hCounter < 539) or (vCounter = 414 and hCounter >= 610 and hCounter < 632) or (vCounter = 415 and hCounter >= 520 and hCounter < 539) or (vCounter = 415 and hCounter >= 611 and hCounter < 633) or (vCounter = 416 and hCounter >= 520 and hCounter < 539) or (vCounter = 416 and hCounter >= 611 and hCounter < 633) or (vCounter = 417 and hCounter >= 520 and hCounter < 539) or (vCounter = 417 and hCounter >= 612 and hCounter < 634) or (vCounter = 418 and hCounter >= 520 and hCounter < 539) or (vCounter = 418 and hCounter >= 612 and hCounter < 634) or (vCounter = 419 and hCounter >= 520 and hCounter < 539) or (vCounter = 419 and hCounter >= 613 and hCounter < 634) or (vCounter = 420 and hCounter >= 520 and hCounter < 539) or (vCounter = 420 and hCounter >= 613 and hCounter < 635) or (vCounter = 421 and hCounter >= 520 and hCounter < 539) or (vCounter = 421 and hCounter >= 614 and hCounter < 635) or (vCounter = 422 and hCounter >= 520 and hCounter < 539) or (vCounter = 422 and hCounter >= 614 and hCounter < 635) or (vCounter = 423 and hCounter >= 520 and hCounter < 539) or (vCounter = 423 and hCounter >= 614 and hCounter < 635) or (vCounter = 424 and hCounter >= 520 and hCounter < 539) or (vCounter = 424 and hCounter >= 615 and hCounter < 636) or (vCounter = 425 and hCounter >= 520 and hCounter < 539) or (vCounter = 425 and hCounter >= 615 and hCounter < 636) or (vCounter = 426 and hCounter >= 520 and hCounter < 539) or (vCounter = 426 and hCounter >= 615 and hCounter < 636) or (vCounter = 427 and hCounter >= 520 and hCounter < 539) or (vCounter = 427 and hCounter >= 616 and hCounter < 637) or (vCounter = 428 and hCounter >= 520 and hCounter < 539) or (vCounter = 428 and hCounter >= 616 and hCounter < 637) or (vCounter = 429 and hCounter >= 520 and hCounter < 539) or (vCounter = 429 and hCounter >= 616 and hCounter < 637) or (vCounter = 430 and hCounter >= 520 and hCounter < 539) or (vCounter = 430 and hCounter >= 617 and hCounter < 637) or (vCounter = 431 and hCounter >= 520 and hCounter < 539) or (vCounter = 431 and hCounter >= 617 and hCounter < 637) or (vCounter = 432 and hCounter >= 520 and hCounter < 539) or (vCounter = 432 and hCounter >= 617 and hCounter < 638) or (vCounter = 433 and hCounter >= 520 and hCounter < 539) or (vCounter = 433 and hCounter >= 617 and hCounter < 638) or (vCounter = 434 and hCounter >= 520 and hCounter < 539) or (vCounter = 434 and hCounter >= 618 and hCounter < 638) or (vCounter = 435 and hCounter >= 520 and hCounter < 539) or (vCounter = 435 and hCounter >= 618 and hCounter < 638) or (vCounter = 436 and hCounter >= 520 and hCounter < 539) or (vCounter = 436 and hCounter >= 618 and hCounter < 638) or (vCounter = 437 and hCounter >= 520 and hCounter < 539) or (vCounter = 437 and hCounter >= 618 and hCounter < 639) or (vCounter = 438 and hCounter >= 520 and hCounter < 539) or (vCounter = 438 and hCounter >= 618 and hCounter < 639) or (vCounter = 439 and hCounter >= 520 and hCounter < 539) or (vCounter = 439 and hCounter >= 619 and hCounter < 639) or (vCounter = 440 and hCounter >= 520 and hCounter < 539) or (vCounter = 440 and hCounter >= 619 and hCounter < 639) or (vCounter = 441 and hCounter >= 520 and hCounter < 539) or (vCounter = 441 and hCounter >= 619 and hCounter < 639) or (vCounter = 442 and hCounter >= 520 and hCounter < 539) or (vCounter = 442 and hCounter >= 619 and hCounter < 639) or (vCounter = 443 and hCounter >= 520 and hCounter < 539) or (vCounter = 443 and hCounter >= 619 and hCounter < 639) or (vCounter = 444 and hCounter >= 520 and hCounter < 539) or (vCounter = 444 and hCounter >= 619 and hCounter < 639) or (vCounter = 445 and hCounter >= 520 and hCounter < 539) or (vCounter = 445 and hCounter >= 619 and hCounter < 639) or (vCounter = 446 and hCounter >= 520 and hCounter < 539) or (vCounter = 446 and hCounter >= 619 and hCounter < 639) or (vCounter = 447 and hCounter >= 520 and hCounter < 539) or (vCounter = 447 and hCounter >= 619 and hCounter < 639) or (vCounter = 448 and hCounter >= 520 and hCounter < 539) or (vCounter = 448 and hCounter >= 619 and hCounter < 639) or (vCounter = 449 and hCounter >= 520 and hCounter < 539) or (vCounter = 449 and hCounter >= 619 and hCounter < 639) or (vCounter = 450 and hCounter >= 520 and hCounter < 539) or (vCounter = 450 and hCounter >= 619 and hCounter < 639) or (vCounter = 451 and hCounter >= 520 and hCounter < 539) or (vCounter = 451 and hCounter >= 620 and hCounter < 639) or (vCounter = 452 and hCounter >= 520 and hCounter < 539) or (vCounter = 452 and hCounter >= 619 and hCounter < 639) or (vCounter = 453 and hCounter >= 520 and hCounter < 539) or (vCounter = 453 and hCounter >= 619 and hCounter < 639) or (vCounter = 454 and hCounter >= 520 and hCounter < 539) or (vCounter = 454 and hCounter >= 619 and hCounter < 639) or (vCounter = 455 and hCounter >= 520 and hCounter < 539) or (vCounter = 455 and hCounter >= 619 and hCounter < 639) or (vCounter = 456 and hCounter >= 520 and hCounter < 539) or (vCounter = 456 and hCounter >= 619 and hCounter < 639) or (vCounter = 457 and hCounter >= 520 and hCounter < 539) or (vCounter = 457 and hCounter >= 619 and hCounter < 639) or (vCounter = 458 and hCounter >= 520 and hCounter < 539) or (vCounter = 458 and hCounter >= 619 and hCounter < 639) or (vCounter = 459 and hCounter >= 520 and hCounter < 539) or (vCounter = 459 and hCounter >= 619 and hCounter < 639) or (vCounter = 460 and hCounter >= 520 and hCounter < 539) or (vCounter = 460 and hCounter >= 619 and hCounter < 639) or (vCounter = 461 and hCounter >= 520 and hCounter < 539) or (vCounter = 461 and hCounter >= 619 and hCounter < 639) or (vCounter = 462 and hCounter >= 520 and hCounter < 539) or (vCounter = 462 and hCounter >= 619 and hCounter < 639) or (vCounter = 463 and hCounter >= 520 and hCounter < 539) or (vCounter = 463 and hCounter >= 619 and hCounter < 639) or (vCounter = 464 and hCounter >= 520 and hCounter < 539) or (vCounter = 464 and hCounter >= 618 and hCounter < 639) or (vCounter = 465 and hCounter >= 520 and hCounter < 539) or (vCounter = 465 and hCounter >= 618 and hCounter < 639) or (vCounter = 466 and hCounter >= 520 and hCounter < 539) or (vCounter = 466 and hCounter >= 618 and hCounter < 638) or (vCounter = 467 and hCounter >= 520 and hCounter < 539) or (vCounter = 467 and hCounter >= 618 and hCounter < 638) or (vCounter = 468 and hCounter >= 520 and hCounter < 539) or (vCounter = 468 and hCounter >= 618 and hCounter < 638) or (vCounter = 469 and hCounter >= 520 and hCounter < 539) or (vCounter = 469 and hCounter >= 617 and hCounter < 638) or (vCounter = 470 and hCounter >= 520 and hCounter < 539) or (vCounter = 470 and hCounter >= 617 and hCounter < 638) or (vCounter = 471 and hCounter >= 520 and hCounter < 539) or (vCounter = 471 and hCounter >= 617 and hCounter < 637) or (vCounter = 472 and hCounter >= 520 and hCounter < 539) or (vCounter = 472 and hCounter >= 617 and hCounter < 637) or (vCounter = 473 and hCounter >= 520 and hCounter < 539) or (vCounter = 473 and hCounter >= 616 and hCounter < 637) or (vCounter = 474 and hCounter >= 520 and hCounter < 539) or (vCounter = 474 and hCounter >= 616 and hCounter < 637) or (vCounter = 475 and hCounter >= 520 and hCounter < 539) or (vCounter = 475 and hCounter >= 616 and hCounter < 637) or (vCounter = 476 and hCounter >= 520 and hCounter < 539) or (vCounter = 476 and hCounter >= 615 and hCounter < 636) or (vCounter = 477 and hCounter >= 520 and hCounter < 539) or (vCounter = 477 and hCounter >= 615 and hCounter < 636) or (vCounter = 478 and hCounter >= 520 and hCounter < 539) or (vCounter = 478 and hCounter >= 615 and hCounter < 636) or (vCounter = 479 and hCounter >= 520 and hCounter < 539) or (vCounter = 479 and hCounter >= 614 and hCounter < 635) or (vCounter = 480 and hCounter >= 520 and hCounter < 539) or (vCounter = 480 and hCounter >= 614 and hCounter < 635) or (vCounter = 481 and hCounter >= 520 and hCounter < 539) or (vCounter = 481 and hCounter >= 614 and hCounter < 635) or (vCounter = 482 and hCounter >= 520 and hCounter < 539) or (vCounter = 482 and hCounter >= 613 and hCounter < 635) or (vCounter = 483 and hCounter >= 520 and hCounter < 539) or (vCounter = 483 and hCounter >= 613 and hCounter < 634) or (vCounter = 484 and hCounter >= 520 and hCounter < 539) or (vCounter = 484 and hCounter >= 612 and hCounter < 634) or (vCounter = 485 and hCounter >= 520 and hCounter < 539) or (vCounter = 485 and hCounter >= 612 and hCounter < 634) or (vCounter = 486 and hCounter >= 520 and hCounter < 539) or (vCounter = 486 and hCounter >= 611 and hCounter < 633) or (vCounter = 487 and hCounter >= 520 and hCounter < 539) or (vCounter = 487 and hCounter >= 611 and hCounter < 633) or (vCounter = 488 and hCounter >= 520 and hCounter < 539) or (vCounter = 488 and hCounter >= 610 and hCounter < 632) or (vCounter = 489 and hCounter >= 520 and hCounter < 539) or (vCounter = 489 and hCounter >= 610 and hCounter < 632) or (vCounter = 490 and hCounter >= 520 and hCounter < 539) or (vCounter = 490 and hCounter >= 609 and hCounter < 632) or (vCounter = 491 and hCounter >= 520 and hCounter < 539) or (vCounter = 491 and hCounter >= 609 and hCounter < 631) or (vCounter = 492 and hCounter >= 520 and hCounter < 539) or (vCounter = 492 and hCounter >= 608 and hCounter < 631) or (vCounter = 493 and hCounter >= 520 and hCounter < 539) or (vCounter = 493 and hCounter >= 608 and hCounter < 630) or (vCounter = 494 and hCounter >= 520 and hCounter < 539) or (vCounter = 494 and hCounter >= 607 and hCounter < 630) or (vCounter = 495 and hCounter >= 520 and hCounter < 539) or (vCounter = 495 and hCounter >= 606 and hCounter < 629) or (vCounter = 496 and hCounter >= 520 and hCounter < 539) or (vCounter = 496 and hCounter >= 606 and hCounter < 629) or (vCounter = 497 and hCounter >= 520 and hCounter < 539) or (vCounter = 497 and hCounter >= 605 and hCounter < 628) or (vCounter = 498 and hCounter >= 520 and hCounter < 539) or (vCounter = 498 and hCounter >= 604 and hCounter < 628) or (vCounter = 499 and hCounter >= 520 and hCounter < 539) or (vCounter = 499 and hCounter >= 604 and hCounter < 627) or (vCounter = 500 and hCounter >= 520 and hCounter < 539) or (vCounter = 500 and hCounter >= 603 and hCounter < 627) or (vCounter = 501 and hCounter >= 520 and hCounter < 539) or (vCounter = 501 and hCounter >= 602 and hCounter < 626) or (vCounter = 502 and hCounter >= 520 and hCounter < 539) or (vCounter = 502 and hCounter >= 601 and hCounter < 626) or (vCounter = 503 and hCounter >= 520 and hCounter < 539) or (vCounter = 503 and hCounter >= 600 and hCounter < 625) or (vCounter = 504 and hCounter >= 520 and hCounter < 539) or (vCounter = 504 and hCounter >= 599 and hCounter < 624) or (vCounter = 505 and hCounter >= 520 and hCounter < 539) or (vCounter = 505 and hCounter >= 599 and hCounter < 624) or (vCounter = 506 and hCounter >= 520 and hCounter < 539) or (vCounter = 506 and hCounter >= 598 and hCounter < 623) or (vCounter = 507 and hCounter >= 520 and hCounter < 539) or (vCounter = 507 and hCounter >= 597 and hCounter < 622) or (vCounter = 508 and hCounter >= 520 and hCounter < 539) or (vCounter = 508 and hCounter >= 596 and hCounter < 622) or (vCounter = 509 and hCounter >= 520 and hCounter < 539) or (vCounter = 509 and hCounter >= 595 and hCounter < 621) or (vCounter = 510 and hCounter >= 520 and hCounter < 539) or (vCounter = 510 and hCounter >= 594 and hCounter < 620) or (vCounter = 511 and hCounter >= 520 and hCounter < 539) or (vCounter = 511 and hCounter >= 592 and hCounter < 619) or (vCounter = 512 and hCounter >= 520 and hCounter < 539) or (vCounter = 512 and hCounter >= 591 and hCounter < 619) or (vCounter = 513 and hCounter >= 520 and hCounter < 539) or (vCounter = 513 and hCounter >= 590 and hCounter < 618) or (vCounter = 514 and hCounter >= 520 and hCounter < 539) or (vCounter = 514 and hCounter >= 589 and hCounter < 617) or (vCounter = 515 and hCounter >= 520 and hCounter < 539) or (vCounter = 515 and hCounter >= 588 and hCounter < 616) or (vCounter = 516 and hCounter >= 520 and hCounter < 539) or (vCounter = 516 and hCounter >= 586 and hCounter < 615) or (vCounter = 517 and hCounter >= 520 and hCounter < 539) or (vCounter = 517 and hCounter >= 585 and hCounter < 615) or (vCounter = 518 and hCounter >= 520 and hCounter < 539) or (vCounter = 518 and hCounter >= 583 and hCounter < 614) or (vCounter = 519 and hCounter >= 520 and hCounter < 539) or (vCounter = 519 and hCounter >= 582 and hCounter < 613) or (vCounter = 520 and hCounter >= 520 and hCounter < 539) or (vCounter = 520 and hCounter >= 580 and hCounter < 612) or (vCounter = 521 and hCounter >= 520 and hCounter < 539) or (vCounter = 521 and hCounter >= 578 and hCounter < 611) or (vCounter = 522 and hCounter >= 520 and hCounter < 539) or (vCounter = 522 and hCounter >= 576 and hCounter < 610) or (vCounter = 523 and hCounter >= 520 and hCounter < 539) or (vCounter = 523 and hCounter >= 574 and hCounter < 609) or (vCounter = 524 and hCounter >= 520 and hCounter < 539) or (vCounter = 524 and hCounter >= 572 and hCounter < 608) or (vCounter = 525 and hCounter >= 520 and hCounter < 539) or (vCounter = 525 and hCounter >= 570 and hCounter < 607) or (vCounter = 526 and hCounter >= 520 and hCounter < 539) or (vCounter = 526 and hCounter >= 567 and hCounter < 606) or (vCounter = 527 and hCounter >= 520 and hCounter < 539) or (vCounter = 527 and hCounter >= 564 and hCounter < 604) or (vCounter = 528 and hCounter >= 520 and hCounter < 539) or (vCounter = 528 and hCounter >= 561 and hCounter < 603) or (vCounter = 529 and hCounter >= 520 and hCounter < 539) or (vCounter = 529 and hCounter >= 557 and hCounter < 602) or (vCounter = 530 and hCounter >= 520 and hCounter < 539) or (vCounter = 530 and hCounter >= 552 and hCounter < 601) or (vCounter = 531 and hCounter >= 520 and hCounter < 539) or (vCounter = 531 and hCounter >= 540 and hCounter < 599) or (vCounter = 532 and hCounter >= 520 and hCounter < 598) or (vCounter = 533 and hCounter >= 520 and hCounter < 597) or (vCounter = 534 and hCounter >= 520 and hCounter < 595) or (vCounter = 535 and hCounter >= 520 and hCounter < 594) or (vCounter = 536 and hCounter >= 520 and hCounter < 592) or (vCounter = 537 and hCounter >= 520 and hCounter < 591) or (vCounter = 538 and hCounter >= 520 and hCounter < 589) or (vCounter = 539 and hCounter >= 520 and hCounter < 587) or (vCounter = 540 and hCounter >= 520 and hCounter < 585) or (vCounter = 541 and hCounter >= 520 and hCounter < 583) or (vCounter = 542 and hCounter >= 520 and hCounter < 581) or (vCounter = 543 and hCounter >= 520 and hCounter < 579) or (vCounter = 544 and hCounter >= 520 and hCounter < 576) or (vCounter = 545 and hCounter >= 520 and hCounter < 574) or (vCounter = 546 and hCounter >= 520 and hCounter < 571) or (vCounter = 547 and hCounter >= 520 and hCounter < 567) or (vCounter = 548 and hCounter >= 520 and hCounter < 564) or (vCounter = 549 and hCounter >= 520 and hCounter < 559) or (vCounter = 550 and hCounter >= 520 and hCounter < 554) then
					--D
					vga_red <= ldispCounter(0);
					vga_green <= ldispCounter(1);
					vga_blue <= ldispCounter(2);
				 elsif (hCounter > 739 and hCounter < 759 and vCounter > 351 and vCounter < 551) or (hCounter > 739 and hCounter < 839 and vCounter> 531 and vCounter < 551) then
					--L
					vga_red <= ldispCounter(0);
					vga_green <= ldispCounter(1);
					vga_blue <= ldispCounter(2);
				 else
					vga_red <= '0';
					vga_green <= '0';
					vga_blue <= '0';
				 end if;
			 end if;
		 else
			vga_red <= '0';
			vga_green <= '0';
			vga_blue <= '0';
		 end if;

		 if vga_shift /= lastShift then
			lastShift <= vga_shift;
			hdispCounter <= hdispCounter + 1;
			vdispCounter <= vdispCounter + 1;
			ldispCounter <= ldispCounter + 1;
		 end if;
		 
		 if vga_state /= lastState then
			state <= state + 1;
			lastState <= vga_state;
		 end if;
		 
		 if state = 3 then
			state <= "00";
		 end if;
		 
      end if;
   end process;
end Behavioral;